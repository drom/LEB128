module pack_i32 ();
endmodule
