module pack_u64 ();

endmodule
