module pack_i64 ();
endmodule
